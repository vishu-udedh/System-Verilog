module AND_GATE(A,B,Y);
input logic A,B;
output logic Y;
assign Y=A&B;
endmodule
